`ifndef _definiciones_vh_
`define _definiciones_vh_
	`define BUS_DAT 8 				//ancho del bus de datos 
	`define BUS_DAT_MSB `BUS_DAT-1 	//ancho del bus de datos MENOS UNO
`endif
